0
0 0 0 0 0 r h 1 B 8 B
0 0 0 0 0 r h 4 B 32 B
0 0 0 0 0 r h 0 B 2 B
0 0 0 0 0 r h 3 B 5 B
4 3 5 7 2 8 2 11 3 4 1 6 0 11 4 2 1 10 3 6 3 12 0 8 2 10 0 9 1 3 4 5 0 5 1 9 2 4
1
